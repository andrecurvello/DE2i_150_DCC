----------------------------------------------------------------------------------
-- Copyright (c) 2014, Luis Ardila
-- E-mail: leardilap@unal.edu.co

-- Revisions: 
-- Date        	Version    	Author    		Description
-- 12/10/2014    	1.0    		Luis Ardila    File created
--
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DE2i_150_DCC_TOP IS 
PORT (
	--	CLOCKS
		CLOCK_50				: IN STD_LOGIC;	
		CLOCK2_50			: IN STD_LOGIC;	
		CLOCK3_50			: IN STD_LOGIC;	

	--	DRAM
		DRAM_ADDR			: OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
		DRAM_BA				: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		DRAM_CAS_N			: OUT STD_LOGIC;
		DRAM_CKE				: OUT STD_LOGIC;
		DRAM_CLK				: OUT STD_LOGIC;
		DRAM_CS_N			: OUT STD_LOGIC;
		DRAM_DQM				: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		DRAM_DQ				: INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
		DRAM_RAS_N			: OUT STD_LOGIC;
		DRAM_WE_N			: OUT STD_LOGIC;

	-- EEP
		EEP_I2C_SCLK		: OUT STD_LOGIC;
		EEP_I2C_SDAT		: INOUT STD_LOGIC;

	-- ENET
		ENET_GTX_CLK		: OUT STD_LOGIC;
		ENET_INT_N			: IN STD_LOGIC;
		ENET_LINK100		: IN STD_LOGIC;
		ENET_MDC				: OUT STD_LOGIC;
		ENET_MDIO			: INOUT STD_LOGIC;
		ENET_RST_N			: OUT STD_LOGIC;
		ENET_RX_CLK			: IN STD_LOGIC;
		ENET_RX_COL			: IN STD_LOGIC;
		ENET_RX_CRS			: IN STD_LOGIC;
		ENET_RX_DATA		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		ENET_RX_DV			: IN STD_LOGIC;
		ENET_RX_ER			: IN STD_LOGIC;
		ENET_TX_CLK			: IN STD_LOGIC;
		ENET_TX_DATA		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		ENET_TX_EN			: OUT STD_LOGIC;
		ENET_TX_ER			: OUT STD_LOGIC;

	-- FAN
		FAN_CTRL				: OUT STD_LOGIC;

	-- FL
		FL_CE_N				: OUT STD_LOGIC;
		FL_OE_N				: OUT STD_LOGIC;
		FL_RESET_N			: OUT STD_LOGIC;
		FL_RY					: IN STD_LOGIC;
		FL_WE_N				: OUT STD_LOGIC;
		FL_WP_N				: OUT STD_LOGIC;

	-- FS
		FS_ADDR				: OUT STD_LOGIC_VECTOR (26 DOWNTO 0);
		FS_DQ					: INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);

	-- GPIO
		GPIO					: INOUT STD_LOGIC_VECTOR (35 DOWNTO 0);

	-- G
		G_SENSOR_INT1		: IN STD_LOGIC;
		G_SENSOR_SCLK		: OUT STD_LOGIC;
		G_SENSOR_SDAT		: INOUT STD_LOGIC;

	-- HEX
		HEX0					: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		HEX1					: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		HEX2					: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		HEX3					: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		HEX4					: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		HEX5					: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		HEX6					: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
		HEX7					: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);

	-- HSMC
		HSMC_CLKIN1			: IN STD_LOGIC; 										--TP1
		HSMC_CLKOUT0		: OUT STD_LOGIC;										--TP2
		HSMC_J1_152			: OUT STD_LOGIC;										--TP5
		
		HSMC_SCL				: OUT STD_LOGIC;
		HSMC_SDA				: INOUT STD_LOGIC;	
		
		HSMC_XT_IN_N		: IN STD_LOGIC;
		HSMC_XT_IN_P		: IN STD_LOGIC;
		
		HSMC_FPGA_CLK_A_N	: OUT STD_LOGIC;
		HSMC_FPGA_CLK_A_P : OUT STD_LOGIC;
		HSMC_FPGA_CLK_B_N	: OUT STD_LOGIC;
		HSMC_FPGA_CLK_B_P : OUT STD_LOGIC;

		HSMC_ADA_D			: IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		HSMC_ADA_OR			: IN STD_LOGIC;
		HSMC_ADA_SPI_CS	: OUT STD_LOGIC;
		HSMC_ADA_OE			: OUT STD_LOGIC;
		HSMC_ADA_DCO		: IN STD_LOGIC;
		
		HSMC_ADB_D			: IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		HSMC_ADB_OR			: IN STD_LOGIC;
		HSMC_ADB_SPI_CS	: OUT STD_LOGIC;
		HSMC_ADB_OE			: OUT STD_LOGIC;
		HSMC_ADB_DCO		: IN STD_LOGIC;
		
		HSMC_DA				: OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
		HSMC_DB				: OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
		
		HSMC_AIC_XCLK		: IN STD_LOGIC;
		HSMC_AIC_LRCOUT	: INOUT STD_LOGIC;
		HSMC_AIC_LRCIN		: INOUT STD_LOGIC;
		HSMC_AIC_DIN		: OUT STD_LOGIC;
		HSMC_AIC_DOUT		: IN STD_LOGIC;
		HSMC_AD_SCLK		: OUT STD_LOGIC;
		HSMC_AD_SDIO		: INOUT STD_LOGIC;
		HSMC_AIC_SPI_CS	: OUT STD_LOGIC;						--low active
		HSMC_AIC_BCLK		: INOUT STD_LOGIC;
		
	-- I2C
		I2C_SCLK				: OUT STD_LOGIC;
		I2C_SDAT				: INOUT STD_LOGIC;

	-- IRDA
		IRDA_RXD				: IN STD_LOGIC;

	-- KEY
		KEY					: IN STD_LOGIC_VECTOR (3 DOWNTO 0);

	-- LCD
		LCD_DATA				: INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		LCD_EN				: OUT STD_LOGIC;
		LCD_ON				: OUT STD_LOGIC;
		LCD_RS				: OUT STD_LOGIC;
		LCD_RW				: OUT STD_LOGIC;

	-- LEDS
		LEDG					: OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
		LEDR					: OUT STD_LOGIC_VECTOR (17 DOWNTO 0);

	-- PCIE
		--PCIE_PERST_N		: IN STD_LOGIC;
		--PCIE_REFCLK_P	: IN STD_LOGIC;
		--PCIE_RX_P			: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		--PCIE_TX_P			: OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		--PCIE_WAKE_N		: OUT STD_LOGIC;

	-- SD
		SD_CLK				: OUT STD_LOGIC;
		SD_CMD				: INOUT STD_LOGIC;
		SD_DAT				: INOUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		SD_WP_N				: IN STD_LOGIC;

	-- SMA
		SMA_CLKIN			: IN STD_LOGIC;
		SMA_CLKOUT        : OUT STD_LOGIC;

	-- SSRAM
		SSRAM0_CE_N       : OUT STD_LOGIC;
		SSRAM1_CE_N       : OUT STD_LOGIC;
		SSRAM_ADSC_N      : OUT STD_LOGIC;
		SSRAM_ADSP_N      : OUT STD_LOGIC;
		SSRAM_ADV_N       : OUT STD_LOGIC;
		SSRAM_BE				: INOUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		SSRAM_CLK			: OUT STD_LOGIC;
		SSRAM_GW_N        : OUT STD_LOGIC;
		SSRAM_OE_N        : OUT STD_LOGIC;
		SSRAM_WE_N        : OUT STD_LOGIC;

	-- SW
		SW						: IN STD_LOGIC_VECTOR (17 DOWNTO 0);

	-- TD
		TD_CLK27				: IN STD_LOGIC;
		TD_DATA				: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		TD_HS					: IN STD_LOGIC;
		TD_RESET_N        : OUT STD_LOGIC;
		TD_VS             : IN STD_LOGIC;

	-- UART
		UART_CTS          : IN STD_LOGIC;
		UART_RTS          : OUT STD_LOGIC;
		UART_RXD          : IN STD_LOGIC;
		UART_TXD          : OUT STD_LOGIC;
		
	-- VGA
		VGA_BLANK_N       : OUT STD_LOGIC;
		VGA_B					: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		VGA_CLK				: OUT STD_LOGIC;
		VGA_G					: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		VGA_HS				: OUT STD_LOGIC;
		VGA_R					: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		VGA_SYNC_N			: OUT STD_LOGIC;
		VGA_VS				: OUT STD_LOGIC
		);
END DE2i_150_DCC_TOP;

ARCHITECTURE DE2i_150_DCC_TOP_ARCH OF DE2i_150_DCC_TOP IS

COMPONENT PLL_1 IS 
PORT (
		inclk0		: IN STD_LOGIC  := '0';
		c0				: OUT STD_LOGIC;
		c1		: OUT STD_LOGIC 
		);
END COMPONENT PLL_1;

COMPONENT HDIG_HEX IS 
PORT (
		HDIG			: IN 	STD_LOGIC_VECTOR (3 DOWNTO 0);
		HEX			: OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
		);
END COMPONENT HDIG_HEX;

COMPONENT AD_SPI_CONTROLLER IS
PORT(
	CLK10					: IN STD_LOGIC;								-- 10 MHz
	RST					: IN STD_LOGIC;
	SPI_ADDRESS			: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	SPI_DATA_IN			: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	SPI_DATA_RW			: IN STD_LOGIC;								--1 READ - 0 WRITE
	SPI_DATA_IN_WEA	: IN STD_LOGIC;
	SPI_DATA_IN_WEB	: IN STD_LOGIC;
	SPI_DATA_OUT		: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	SPI_DATA_OUT_WEA	: OUT STD_LOGIC;
	SPI_DATA_OUT_WEB	: OUT STD_LOGIC;
	SPI_BUSY				: OUT STD_LOGIC;
	-- ADCs SPI INTERFACE
	AD_SCLK				: OUT STD_LOGIC;
	AD_SDIO				: INOUT STD_LOGIC;
	ADA_SPI_CS_n		: OUT STD_LOGIC;
	ADB_SPI_CS_n		: OUT STD_LOGIC
	);
END COMPONENT AD_SPI_CONTROLLER;

COMPONENT LCD16x2 IS 
GENERIC (
  CLK_PERIOD_NS : POSITIVE := 20);    -- 50MHz   --POSITIVE is INTEGER but from 1 to 2147483647
PORT (	
  CLK            : IN STD_LOGIC;
  RST            : IN STD_LOGIC;
	ADA_DATA_IN    : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
	ADA_DATA_EN    : IN STD_LOGIC;
	ADB_DATA_IN			 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
	ADB_DATA_EN    : IN STD_LOGIC;    
	--LCD INTERFACE
	LCD_DATA       : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
	LCD_EN				     : OUT STD_LOGIC;
	LCD_ON				     : OUT STD_LOGIC;
	LCD_RS				     : OUT STD_LOGIC;
	LCD_RW				     : OUT STD_LOGIC
	);
END COMPONENT LCD16x2;

-- SIGNALs FOR OUTSIDE
SIGNAL	RST			:	STD_LOGIC; 	
SIGNAL	SUB			:	STD_LOGIC; 	
SIGNAL	ADD         :	STD_LOGIC; 	
SIGNAL	SEG_0		:	STD_LOGIC_VECTOR (6 DOWNTO 0); --Seven Segments ¨HEX0¨ 

SIGNAL sCLK10 				: STD_LOGIC := '0';
SIGNAL sCLK5k 				: STD_LOGIC := '0';
SIGNAL sADD					: 	STD_LOGIC := '0';
SIGNAL sSUB					: 	STD_LOGIC := '0';
SIGNAL sHDIG				:	STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
SIGNAL sHEX0				:	STD_LOGIC_VECTOR (6 DOWNTO 0) := (OTHERS => '0');
SIGNAL sHEX2				:	STD_LOGIC_VECTOR (6 DOWNTO 0) := (OTHERS => '0');
SIGNAL sHEX3				:	STD_LOGIC_VECTOR (6 DOWNTO 0) := (OTHERS => '0');
SIGNAL sHEX4				:	STD_LOGIC_VECTOR (6 DOWNTO 0) := (OTHERS => '0');
SIGNAL sHEX5				:	STD_LOGIC_VECTOR (6 DOWNTO 0) := (OTHERS => '0');
SIGNAL sHEX6				:	STD_LOGIC_VECTOR (6 DOWNTO 0) := (OTHERS => '0');
SIGNAL sHEX7				:	STD_LOGIC_VECTOR (6 DOWNTO 0) := (OTHERS => '0');

SIGNAL sSPI_DATA_OUT  		: STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
SIGNAL sSPI_DATA_IN_WEA		: STD_LOGIC := '0';
SIGNAL sSPI_DATA_OUT_WEA	: STD_LOGIC := '0';
SIGNAL sSPI_DATA_OUT_WEB	: STD_LOGIC := '0';
SIGNAL sSPI_BUSY				: STD_LOGIC := '0';

SIGNAL sSPI_CNT  				: INTEGER RANGE 0 to 65500 := 0;

BEGIN 

PLL_1_inst : PLL_1 
PORT MAP (
		inclk0	=> CLOCK_50,
		c0	 		=> sCLK10,
		c1			=> sCLK5k
		);

HEX0_Inst : HDIG_HEX 
PORT MAP (
		HDIG	=> sHDIG,
		HEX	=> sHEX0
		);
		
AD_SPI_CONTROLLER_inst : AD_SPI_CONTROLLER
PORT MAP (
	CLK10						=> sCLK10,
	RST						=> RST,
	SPI_ADDRESS				=> SW(15 DOWNTO 8),
	SPI_DATA_IN				=> SW(7 DOWNTO 0),
	SPI_DATA_RW				=> SW(17),							--1 READ - 0 WRITE
	SPI_DATA_IN_WEA	   => sSPI_DATA_IN_WEA,
	SPI_DATA_IN_WEB	   => '0',
	SPI_DATA_OUT			=> sSPI_DATA_OUT,
	SPI_DATA_OUT_WEA		=> sSPI_DATA_OUT_WEA,
	SPI_DATA_OUT_WEB		=> sSPI_DATA_OUT_WEB,
	SPI_BUSY					=> sSPI_BUSY,
	-- ADCs SPI INTERFACE
	AD_SCLK					=> HSMC_AD_SCLK,	
	AD_SDIO					=> HSMC_AD_SDIO,			
	ADA_SPI_CS_n			=> HSMC_ADA_SPI_CS,
	ADB_SPI_CS_n			=> HSMC_ADB_SPI_CS
	);
	
LCD16x2_INST : LCD16x2
GENERIC MAP(
	CLK_PERIOD_NS => 100)    -- 10MHz   --POSITIVE is INTEGER but from 1 to 2147483647
PORT MAP(	
	CLK            => sCLK10,
	RST            => RST,
	ADA_DATA_IN    => sSPI_DATA_OUT,
	ADA_DATA_EN    => sSPI_DATA_OUT_WEA,
	ADB_DATA_IN		=> sSPI_DATA_OUT,
	ADB_DATA_EN    => sSPI_DATA_OUT_WEB,   
	--LCD INTERFACE
	LCD_DATA       => LCD_DATA,
	LCD_EN			=> LCD_EN,
	LCD_ON			=> LCD_ON,
	LCD_RS			=> LCD_RS,
	LCD_RW			=> LCD_RW
	);

HEX2_Inst : HDIG_HEX 
PORT MAP (
		HDIG	=> sSPI_DATA_OUT(3 DOWNTO 0),
		HEX	=> sHEX2
		);

HEX3_Inst : HDIG_HEX 
PORT MAP (
		HDIG	=> sSPI_DATA_OUT(7 DOWNTO 4),
		HEX	=> sHEX3
		);
		
HEX4_Inst : HDIG_HEX 
PORT MAP (
		HDIG	=> SW(3 DOWNTO 0),
		HEX	=> sHEX4
		);

HEX5_Inst : HDIG_HEX 
PORT MAP (
		HDIG	=> SW(7 DOWNTO 4),
		HEX	=> sHEX5
		);
		
HEX6_Inst : HDIG_HEX 
PORT MAP (
		HDIG	=> SW(11 DOWNTO 8),
		HEX	=> sHEX6
		);

HEX7_Inst : HDIG_HEX 
PORT MAP (
		HDIG	=> SW(15 DOWNTO 12),
		HEX	=> sHEX7
		);

AD_SPI_PROCESS : PROCESS (sCLK10, RST) IS
BEGIN
	IF RST = '1' THEN
		sSPI_DATA_IN_WEA <= '0';
	ELSIF rising_edge(sCLK10) AND sSPI_BUSY = '0' THEN
		sSPI_DATA_IN_WEA <= '0';
		IF KEY(3) = '0' THEN
			IF sSPI_CNT > 65000 THEN
				sSPI_DATA_IN_WEA <= '1';
				sSPI_CNT <= 0;
			ELSE 
				sSPI_DATA_IN_WEA <= '0';
				sSPI_CNT <= sSPI_CNT + 1;
			END IF;
		END IF;
	END IF;
	
END PROCESS AD_SPI_PROCESS;

COUNTER: PROCESS (sCLK10, RST) IS
BEGIN

	IF RST = '1' THEN
		sHDIG <= (OTHERS => '0');
	ELSIF rising_edge(sCLK10) THEN
		sADD <= ADD;
		sSUB <= SUB;
		IF (sADD = '1') AND (ADD = '0')  AND (SUB = '1') THEN							--add
			sHDIG <= STD_LOGIC_VECTOR(UNSIGNED(sHDIG) + 1);
		ELSIF (sSUB = '1') AND (SUB = '0') AND (ADD = '1') THEN						--subtract
			sHDIG <= STD_LOGIC_VECTOR(UNSIGNED(sHDIG) - 1);
		ELSE
			sHDIG <= sHDIG;													--keep value
		END IF;
	END IF;
END PROCESS COUNTER;

RST		<= not KEY(2);
SUB		<= KEY(1);
ADD		<= KEY(0); 

LEDR		<= SW;
LEDG 		<= b"00" & sHEX0;

HEX0 		<= sHEX0;
HEX1		<= (OTHERS => '1');
HEX2		<= sHEX2;
HEX3		<= sHEX3;
HEX4		<= sHEX4;
HEX5		<= sHEX5;
HEX6		<= sHEX6;
HEX7		<= sHEX7;

--Turn fan off
FAN_CTRL <= '0';

END DE2i_150_DCC_TOP_ARCH;